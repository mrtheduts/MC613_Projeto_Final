package common is

	type estado_t is (subindo, descendo);

end common;

package body common is
--nada
end common;